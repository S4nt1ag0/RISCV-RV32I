//componente para gerar imediato de 32 bits
//componente para gerar os sinais de controle
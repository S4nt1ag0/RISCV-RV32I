//------------------------------------------------------------------------------
// Definitions and macros for RISCV agent
//------------------------------------------------------------------------------
// This file contains definitions and macros used by the RISCV agent.
//
// Author: Gustavo Santiago
// Date  : June 2025
//------------------------------------------------------------------------------

`ifndef RISCV_DEFINES
`define RISCV_DEFINES

  `define RISCV_WIDTH 4 
  `define NO_OF_TRANSACTIONS 1000

`endif

//componente para gerar instruction decode